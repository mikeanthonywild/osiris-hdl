/* 
 * top.v
 *
 * Author: Mike Wild <m.a.wild@se12.qmul.ac.uk>
 * Date: 14th October 2015
 *
 * This is the top-level module for the OV7670 camera module, comprising of 
 * miniSpartan 6+ development board and OV7670 image sensor.
 */

